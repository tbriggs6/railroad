** Profile: "SCHEMATIC1-bias"  [ C:\orcad_projects\Railroad\raillroad-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\tbriggs\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "C:\orcad\libraries\pspice\TPS2051B_PSPICE_TRANS\tps2051b_sot235.lib" 
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10m 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
